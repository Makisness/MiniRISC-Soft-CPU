module main (
    
);
    
endmodule